module vga_controller(iRST_n,
                      iVGA_CLK,
                      oBLANK_n,
                      oHS,
                      oVS,
                      b_data,
                      g_data,
                      r_data,write_clock,
               write_addr,
               write_data,
               wren_signal);
input iRST_n;
input iVGA_CLK;
input wren_signal;
input write_clock;
output reg oBLANK_n;
output reg oHS;
output reg oVS;
input [18:0] write_addr;
input [23:0] write_data;
output [7:0] b_data;
output [7:0] g_data;  
output [7:0] r_data;                        
///////// ////                     
reg [18:0] ADDR;
reg [23:0] bgr_data;
wire VGA_CLK_n;
wire [7:0] index;
wire [23:0] bgr_data_raw;
wire cBLANK_n,cHS,cVS,rst;
////
assign rst = ~iRST_n;
video_sync_generator LTM_ins (.vga_clk(iVGA_CLK),
                              .reset(rst),
                              .blank_n(cBLANK_n),
                              .HS(cHS),
                              .VS(cVS));
////
////Addresss generator
always@(posedge iVGA_CLK,negedge iRST_n)
begin
  if (!iRST_n)
     ADDR<=19'd0;
  else if (cHS==1'b0 && cVS==1'b0)
     ADDR<=19'd0;
  else if (cBLANK_n==1'b1)
     ADDR<=ADDR+1;
end
//////////////////////////
//////INDEX addr.
assign VGA_CLK_n = ~iVGA_CLK;
img_data_final img_data_memory(
  .address_a(ADDR),
  .address_b(write_addr),
  .clock_a(VGA_CLK_n),
  .clock_b(write_clock),
  .data_b(write_data),
  .wren_b(wren_signal),
  .q_a(index));
  
//img_data  img_data_inst (
//  .address ( ADDR ),
//  .clock ( VGA_CLK_n ),
//  .q ( index )
//  );
  
//////Color table output
img_index img_index_inst (
  .address ( index ),
  .clock ( iVGA_CLK ),
  .q ( bgr_data_raw)
  );  
//////
//////latch valid data at falling edge;
always@(posedge VGA_CLK_n) bgr_data <= bgr_data_raw;
assign b_data = bgr_data[23:16];
assign g_data = bgr_data[15:8];
assign r_data = bgr_data[7:0];
///////////////////
//////Delay the iHD, iVD,iDEN for one clock cycle;
always@(negedge iVGA_CLK)
begin
  oHS<=cHS;
  oVS<=cVS;
  oBLANK_n<=cBLANK_n;
end

endmodule
  
















