module mult_stall_logic()


endmodule