library verilog;
use verilog.vl_types.all;
entity testbench_jw is
end testbench_jw;
