library verilog;
use verilog.vl_types.all;
entity decoder5to32_vlg_vec_tst is
end decoder5to32_vlg_vec_tst;
