library verilog;
use verilog.vl_types.all;
entity regfile_tb is
end regfile_tb;
