library verilog;
use verilog.vl_types.all;
entity booth_decoder_vlg_vec_tst is
end booth_decoder_vlg_vec_tst;
