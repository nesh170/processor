module control_writeback(instruction,write_reg_number,jal_signal,lw_signal,wren_signal);
	input[31:0] instruction;
	output[4:0] write_reg_number;
	output jal_signal,lw_signal,wren_signal;
	
	
	
	
endmodule