library verilog;
use verilog.vl_types.all;
entity shift_right_arithmetic_vlg_vec_tst is
end shift_right_arithmetic_vlg_vec_tst;
