library verilog;
use verilog.vl_types.all;
entity subtractor_32bit_vlg_vec_tst is
end subtractor_32bit_vlg_vec_tst;
