library verilog;
use verilog.vl_types.all;
entity sl290_hw1_vlg_vec_tst is
end sl290_hw1_vlg_vec_tst;
