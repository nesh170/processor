library verilog;
use verilog.vl_types.all;
entity carry_select_Adder_vlg_vec_tst is
end carry_select_Adder_vlg_vec_tst;
