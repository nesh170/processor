library verilog;
use verilog.vl_types.all;
entity shift_left_logical_vlg_vec_tst is
end shift_left_logical_vlg_vec_tst;
